-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Monday, April 27, 2020 13:53:22 Hora de verano romance

